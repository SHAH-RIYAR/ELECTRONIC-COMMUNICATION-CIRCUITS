CircuitMaker Text
5.6
Probes: 3
V1_1
Transient Analysis
0 165 137 255
V2_1
Transient Analysis
1 177 271 16711680
C3_2
Transient Analysis
2 601 133 32768
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.389325 0.500000
344 176 1532 424
9961490 0
0
6 Title:
5 Name:
0
0
0
29
7 Ground~
168 372 344 0 1 3
0 2
0
0 0 53344 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5130 0 0
2
45641.4 0
0
8 Battery~
219 374 306 0 2 5
0 2 4
0
0 0 864 180
2 8V
14 -2 28 6
2 V4
15 -12 29 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
391 0 0
2
45641.4 1
0
13 Var Resistor~
219 274 270 0 3 7
0 5 4 6
0
0 0 832 180
7 50k 50%
-25 -22 24 -14
3 R13
-11 -32 10 -24
0
0
32 %DA %1 %2 25000
%DB %2 %3 25000
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
82 0 0 0 1 0 0 0
1 R
3124 0 0
2
45641.4 2
0
7 Ground~
168 351 256 0 1 3
0 2
0
0 0 53344 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3421 0 0
2
45641.4 3
0
7 Ground~
168 558 314 0 1 3
0 2
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8157 0 0
2
45641.4 4
0
10 Capacitor~
219 606 162 0 2 5
0 10 8
0
0 0 832 90
5 0.1uF
11 0 46 8
2 C3
22 -10 36 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5572 0 0
2
45641.4 5
0
7 Ground~
168 598 28 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8901 0 0
2
45641.4 6
0
8 Battery~
219 543 29 0 2 5
0 11 2
0
0 0 864 180
3 12V
11 -2 32 6
2 V3
15 -12 29 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7361 0 0
2
45641.4 7
0
7 Ground~
168 287 92 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4747 0 0
2
45641.4 8
0
7 Ground~
168 211 72 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
972 0 0
2
45641.4 9
0
10 Capacitor~
219 287 64 0 2 5
0 2 13
0
0 0 832 90
5 0.1uF
11 0 46 8
2 C2
22 -10 36 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3472 0 0
2
45641.4 10
0
10 Capacitor~
219 190 136 0 2 5
0 17 16
0
0 0 832 0
5 0.1uF
-18 -18 17 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9998 0 0
2
45641.4 11
0
6 MC1496
219 433 197 0 10 21
0 15 13 16 7 3 4 9 12 8
14
0
0 0 4800 0
6 MC1496
-21 -42 21 -34
2 U1
-7 -43 7 -35
0
0
36 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %10 %S
0
0
5 DIP14
21

0 2 8 10 1 4 14 5 12 6
3 2 8 10 1 4 14 5 12 6
3 0
88 0 0 0 1 0 0 0
1 U
3536 0 0
2
45641.4 12
0
7 Ground~
168 197 313 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
45641.4 13
0
7 Ground~
168 159 162 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3835 0 0
2
45641.4 14
0
11 Signal Gen~
195 123 277 0 64 64
0 7 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1167867904 0 1050253722
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 5000 0 0.3 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
11 -300m/300mV
-39 -30 38 -22
2 V2
-7 -40 7 -32
0
0
39 %D %1 %2 DC 0 SIN(0 300m 5k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3670 0 0
2
45641.4 15
0
11 Signal Gen~
195 110 140 0 19 64
0 17 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1195593728 0 1058642330
20
1 50000 0 0.6 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
11 -600m/600mV
-39 -30 38 -22
2 V1
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(0 600m 50k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
5616 0 0
2
45641.4 16
0
9 Resistor~
219 227 231 0 2 5
0 6 7
0
0 0 864 90
3 750
5 0 26 8
3 R12
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9323 0 0
2
45641.4 17
0
9 Resistor~
219 296 218 0 2 5
0 5 3
0
0 0 864 90
3 750
5 0 26 8
3 R11
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
317 0 0
2
45641.4 18
0
9 Resistor~
219 333 223 0 3 5
0 2 7 -1
0
0 0 864 90
2 51
8 0 22 8
3 R10
7 -11 28 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3108 0 0
2
45641.4 19
0
9 Resistor~
219 368 222 0 3 5
0 2 3 -1
0
0 0 864 90
2 51
8 0 22 8
2 R9
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4299 0 0
2
45641.4 20
0
9 Resistor~
219 537 225 0 3 5
0 2 9 -1
0
0 0 864 90
4 6.8k
8 0 36 8
2 R8
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9672 0 0
2
45641.4 21
0
9 Resistor~
219 606 220 0 3 5
0 2 10 -1
0
0 0 864 90
4 6.8k
8 0 36 8
2 R7
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7876 0 0
2
45641.4 22
0
9 Resistor~
219 584 78 0 2 5
0 12 11
0
0 0 864 90
4 3.9k
14 3 42 11
2 R6
23 -10 37 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6369 0 0
2
45641.4 23
0
9 Resistor~
219 517 86 0 2 5
0 8 11
0
0 0 864 90
4 3.9k
4 1 32 9
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9172 0 0
2
45641.4 24
0
9 Resistor~
219 429 49 0 2 5
0 13 11
0
0 0 864 0
4 1000
-14 -14 14 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7100 0 0
2
45641.4 25
0
9 Resistor~
219 245 49 0 3 5
0 2 13 -1
0
0 0 864 0
4 1000
-14 -14 14 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3820 0 0
2
45641.4 26
0
9 Resistor~
219 431 83 0 2 5
0 15 14
0
0 0 864 0
4 1000
-14 -14 14 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7678 0 0
2
45641.4 27
0
9 Resistor~
219 335 121 0 2 5
0 16 13
0
0 0 864 0
2 51
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
961 0 0
2
45641.4 28
0
36
1 0 2 0 0 4096 0 4 0 0 11 3
351 250
351 240
349 240
2 0 3 0 0 4096 0 21 0 0 8 2
368 204
368 160
2 0 4 0 0 4096 0 2 0 0 5 2
372 291
372 274
1 1 2 0 0 12288 0 2 1 0 0 4
372 315
372 314
372 314
372 338
2 6 4 0 0 4224 0 3 13 0 0 4
276 274
482 274
482 215
465 215
1 1 5 0 0 4224 0 19 3 0 0 3
296 236
296 262
292 262
1 3 6 0 0 8320 0 18 3 0 0 3
227 249
227 262
256 262
5 2 3 0 0 16512 0 13 19 0 0 6
401 215
401 163
368 163
368 160
296 160
296 200
2 0 7 0 0 8192 0 18 0 0 12 3
227 213
227 197
199 197
2 0 7 0 0 4096 0 20 0 0 12 2
333 205
333 151
1 1 2 0 0 8192 0 20 21 0 0 3
333 241
333 240
368 240
1 4 7 0 0 12416 0 16 13 0 0 7
154 272
199 272
199 151
333 151
333 190
401 190
401 206
1 0 2 0 0 8192 0 5 0 0 16 3
558 308
557 308
557 262
0 2 8 0 0 4096 0 0 6 22 0 3
517 133
606 133
606 153
7 2 9 0 0 4224 0 13 22 0 0 3
465 206
537 206
537 207
1 1 2 0 0 8320 0 22 23 0 0 4
537 243
537 262
606 262
606 238
1 2 10 0 0 4224 0 6 23 0 0 2
606 171
606 202
2 1 2 0 0 0 0 8 7 0 0 4
541 14
541 9
598 9
598 22
1 0 11 0 0 4096 0 8 0 0 20 2
541 38
541 49
2 0 11 0 0 8320 0 24 0 0 23 3
584 60
584 49
503 49
8 1 12 0 0 4224 0 13 24 0 0 3
465 197
584 197
584 96
1 9 8 0 0 4224 0 25 13 0 0 4
517 104
517 245
465 245
465 188
2 2 11 0 0 0 0 26 25 0 0 3
447 49
517 49
517 68
1 0 13 0 0 4096 0 26 0 0 26 2
411 49
366 49
2 0 13 0 0 0 0 11 0 0 26 2
287 55
287 49
2 0 13 0 0 4224 0 27 0 0 31 3
263 49
367 49
367 121
1 1 2 0 0 0 0 11 9 0 0 2
287 73
287 86
1 1 2 0 0 0 0 27 10 0 0 3
227 49
211 49
211 66
10 2 14 0 0 8320 0 13 28 0 0 4
465 179
470 179
470 83
449 83
1 1 15 0 0 8320 0 28 13 0 0 4
413 83
395 83
395 179
401 179
2 2 13 0 0 0 0 29 13 0 0 4
353 121
389 121
389 188
401 188
1 0 16 0 0 8192 0 29 0 0 33 3
317 121
305 121
305 135
2 3 16 0 0 4224 0 12 13 0 0 6
199 136
305 136
305 135
384 135
384 197
401 197
1 1 17 0 0 4224 0 12 17 0 0 4
181 136
156 136
156 135
141 135
2 1 2 0 0 0 0 16 14 0 0 3
154 282
197 282
197 307
2 1 2 0 0 0 0 17 15 0 0 3
141 145
159 145
159 156
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
14 49 205 73
21 54 197 70
22 NAME: SHAHRIYAR SHAHID
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
37 25 132 49
44 30 124 46
10 MODULATION
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.001 2e-06 2e-06
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
