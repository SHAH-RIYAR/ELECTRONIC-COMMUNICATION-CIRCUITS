CircuitMaker Text
5.6
Probes: 3
V1_1
Transient Analysis
0 139 121 255
V2_1
Transient Analysis
1 125 289 16711680
C3_2
Transient Analysis
2 712 113 32768
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 80 30 150 10
176 80 1364 390
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 2 0.500000 0.500000
344 176 1532 494
9961490 0
0
6 Title:
5 Name:
0
0
0
35
7 Ground~
168 300 368 0 1 3
0 2
0
0 0 53360 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5130 0 0
2
5.90151e-315 0
0
8 Battery~
219 302 320 0 2 5
0 2 7
0
0 0 880 180
2 8V
14 -2 28 6
2 V4
15 -12 29 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
391 0 0
2
5.90151e-315 5.26354e-315
0
7 Ground~
168 314 266 0 1 3
0 2
0
0 0 53360 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3124 0 0
2
5.90151e-315 5.30499e-315
0
13 Var Resistor~
219 235 273 0 3 7
0 9 7 10
0
0 0 848 180
7 50k 50%
-25 -22 24 -14
3 R13
-11 -32 10 -24
0
0
32 %DA %1 %2 25000
%DB %2 %3 25000
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
82 0 0 0 1 0 0 0
1 R
3421 0 0
2
5.90151e-315 5.32571e-315
0
7 Ground~
168 443 275 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8157 0 0
2
5.90151e-315 5.34643e-315
0
10 Capacitor~
219 472 149 0 2 5
0 12 13
0
0 0 848 90
5 0.1uF
4 0 39 8
2 C6
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 22
67 0 0 0 1 0 0 0
1 C
5572 0 0
2
5.90151e-315 5.3568e-315
0
7 Ground~
168 566 298 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8901 0 0
2
5.90151e-315 5.36716e-315
0
10 Capacitor~
219 525 178 0 2 5
0 2 4
0
0 0 848 90
7 0.001uF
10 5 59 13
2 C5
26 -8 40 0
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 62
67 0 0 0 1 0 0 0
1 C
7361 0 0
2
5.90151e-315 5.37752e-315
0
10 Capacitor~
219 600 181 0 2 5
0 2 3
0
0 0 848 90
7 0.001uF
6 8 55 16
2 C4
21 -4 35 4
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 250
67 0 0 0 1 0 0 0
1 C
4747 0 0
2
5.90151e-315 5.38788e-315
0
10 Capacitor~
219 665 113 0 2 5
0 3 14
0
0 0 848 0
6 0.01uF
-21 -18 21 -10
2 C3
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 250
67 0 0 0 1 0 0 0
1 C
972 0 0
2
5.90151e-315 5.39306e-315
0
7 Ground~
168 564 27 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3472 0 0
2
5.90151e-315 5.39824e-315
0
8 Battery~
219 440 32 0 2 5
0 15 2
0
0 0 880 180
3 12V
11 -2 32 6
2 V3
15 -12 29 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
9998 0 0
2
5.90151e-315 5.40342e-315
0
7 Ground~
168 229 76 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3536 0 0
2
5.90151e-315 5.4086e-315
0
7 Ground~
168 82 59 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
5.90151e-315 5.41378e-315
0
10 Capacitor~
219 230 51 0 2 5
0 2 17
0
0 0 848 90
5 0.1uF
9 0 44 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 62
67 0 0 0 1 0 0 0
1 C
3835 0 0
2
5.90151e-315 5.41896e-315
0
6 MC1496
219 347 151 0 10 21
0 19 17 16 5 8 7 11 4 13
18
0
0 0 4816 0
6 MC1496
-21 -42 21 -34
2 U1
-7 -43 7 -35
0
0
36 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %10 %S
0
0
5 DIP14
21

0 2 8 10 1 4 14 5 12 6
3 2 8 10 1 4 14 5 12 6
3 0
88 0 0 0 1 0 0 0
1 U
3670 0 0
2
5.90151e-315 5.42414e-315
0
10 Capacitor~
219 174 121 0 2 5
0 6 16
0
0 0 848 0
5 0.1uF
-18 -18 17 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 62
67 0 0 0 1 0 0 0
1 C
5616 0 0
2
5.90151e-315 5.42933e-315
0
7 Ground~
168 190 341 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9323 0 0
2
5.90151e-315 5.43192e-315
0
7 Ground~
168 150 211 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
317 0 0
2
5.90151e-315 5.43451e-315
0
11 Signal Gen~
195 78 294 0 64 64
0 5 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1203982336 0 1063675494
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 100000 0 0.9 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
11 -900m/900mV
-39 -30 38 -22
2 V2
-7 -40 7 -32
0
0
41 %D %1 %2 DC 0 SIN(0 900m 100k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3108 0 0
2
5.90151e-315 5.4371e-315
0
11 Signal Gen~
195 76 192 0 19 64
0 6 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 0 1203982336 0 1008981770
20
0 100000 0 0.01 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -10m/10mV
-31 -30 32 -22
2 V1
-7 -40 7 -32
0
0
33 %D %1 %2 DC 0 SIN(0 10m 100k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
4299 0 0
2
5.90151e-315 5.43969e-315
0
9 Resistor~
219 297 213 0 3 5
0 2 5 -1
0
0 0 880 90
2 51
11 0 25 8
3 R15
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9672 0 0
2
5.90151e-315 5.44228e-315
0
9 Resistor~
219 330 213 0 3 5
0 2 8 -1
0
0 0 880 90
2 51
11 0 25 8
3 R14
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 70
82 0 0 0 1 0 0 0
1 R
7876 0 0
2
5.90151e-315 5.44487e-315
0
9 Resistor~
219 258 212 0 2 5
0 9 8
0
0 0 880 90
3 750
8 0 29 8
3 R12
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6369 0 0
2
5.90151e-315 5.44746e-315
0
9 Resistor~
219 211 214 0 2 5
0 10 5
0
0 0 880 90
3 750
8 0 29 8
3 R11
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 104226052
82 0 0 0 1 0 0 0
1 R
9172 0 0
2
5.90151e-315 5.45005e-315
0
9 Resistor~
219 414 206 0 3 5
0 2 11 -1
0
0 0 880 90
4 6.8k
4 0 32 8
3 R10
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 62
82 0 0 0 1 0 0 0
1 R
7100 0 0
2
5.90151e-315 5.45264e-315
0
9 Resistor~
219 472 206 0 3 5
0 2 12 -1
0
0 0 880 90
4 6.8k
2 0 30 8
2 R9
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 18
82 0 0 0 1 0 0 0
1 R
3820 0 0
2
5.90151e-315 5.45523e-315
0
9 Resistor~
219 719 179 0 3 5
0 2 14 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R8
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 250
82 0 0 0 1 0 0 0
1 R
7678 0 0
2
5.90151e-315 5.45782e-315
0
9 Resistor~
219 551 113 0 2 5
0 4 3
0
0 0 880 0
4 1000
-14 -14 14 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 250
82 0 0 0 1 0 0 0
1 R
961 0 0
2
5.90151e-315 5.46041e-315
0
9 Resistor~
219 449 82 0 2 5
0 4 15
0
0 0 880 90
4 3.9k
4 1 32 9
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3178 0 0
2
5.90151e-315 5.463e-315
0
9 Resistor~
219 175 32 0 3 5
0 2 17 -1
0
0 0 880 0
4 1000
-14 -14 14 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 18
82 0 0 0 1 0 0 0
1 R
3409 0 0
2
5.90151e-315 5.46559e-315
0
9 Resistor~
219 404 83 0 2 5
0 13 15
0
0 0 880 90
4 3.9k
1 0 29 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 18
82 0 0 0 1 0 0 0
1 R
3951 0 0
2
5.90151e-315 5.46818e-315
0
9 Resistor~
219 322 33 0 2 5
0 17 15
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 18
82 0 0 0 1 0 0 0
1 R
8885 0 0
2
5.90151e-315 5.47077e-315
0
9 Resistor~
219 328 75 0 2 5
0 19 18
0
0 0 880 0
4 1000
-14 -14 14 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 62
82 0 0 0 1 0 0 0
1 R
3780 0 0
2
5.90151e-315 5.47207e-315
0
9 Resistor~
219 236 114 0 2 5
0 16 17
0
0 0 880 0
2 51
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 18
82 0 0 0 1 0 0 0
1 R
9265 0 0
2
5.90151e-315 5.47336e-315
0
44
0 1 2 0 0 4096 0 0 5 21 0 2
443 231
443 269
0 1 2 0 0 0 0 0 3 12 0 2
314 245
314 260
1 0 2 0 0 4096 0 7 0 0 24 2
566 292
566 238
0 1 2 0 0 8192 0 0 28 24 0 4
598 238
598 239
719 239
719 197
0 2 3 0 0 4096 0 0 9 7 0 2
600 113
600 172
0 2 4 0 0 4096 0 0 8 26 0 2
525 113
525 169
2 1 3 0 0 4224 0 29 10 0 0 2
569 113
656 113
1 0 5 0 0 8192 0 20 0 0 19 3
109 289
176 289
176 196
1 1 6 0 0 8320 0 17 21 0 0 3
165 121
107 121
107 187
2 0 7 0 0 4096 0 2 0 0 15 4
300 305
300 297
299 297
299 294
1 1 2 0 0 0 0 2 1 0 0 2
300 329
300 362
1 1 2 0 0 0 0 22 23 0 0 4
297 231
297 245
330 245
330 231
2 0 8 0 0 8192 0 23 0 0 18 4
330 195
330 178
287 178
287 143
2 4 5 0 0 0 0 22 16 0 0 6
297 195
278 195
278 134
278 134
278 160
315 160
2 6 7 0 0 8320 0 4 16 0 0 5
237 277
237 294
382 294
382 169
379 169
1 1 9 0 0 8320 0 4 24 0 0 3
253 265
258 265
258 230
1 3 10 0 0 4224 0 25 4 0 0 3
211 232
211 265
217 265
2 5 8 0 0 4224 0 24 16 0 0 5
258 194
258 143
287 143
287 169
315 169
2 0 5 0 0 12416 0 25 0 0 14 4
211 196
176 196
176 134
278 134
7 2 11 0 0 4224 0 16 26 0 0 3
379 160
414 160
414 188
1 1 2 0 0 0 0 26 27 0 0 4
414 224
414 231
472 231
472 224
1 2 12 0 0 4224 0 6 27 0 0 2
472 158
472 188
2 0 13 0 0 4224 0 6 0 0 37 4
472 140
421 140
421 116
402 116
1 1 2 0 0 0 0 8 9 0 0 4
525 187
525 238
600 238
600 190
2 2 14 0 0 8320 0 10 28 0 0 3
674 113
719 113
719 161
1 0 4 0 0 0 0 29 0 0 30 4
533 113
479 113
479 115
443 115
1 0 15 0 0 4096 0 12 0 0 29 2
438 41
438 52
2 1 2 0 0 4224 0 12 11 0 0 3
438 17
564 17
564 21
0 2 15 0 0 4096 0 0 30 38 0 3
403 52
449 52
449 64
8 1 4 0 0 4224 0 16 30 0 0 5
379 151
443 151
443 115
449 115
449 100
1 0 16 0 0 4096 0 35 0 0 42 3
218 114
211 114
211 121
0 0 17 0 0 4096 0 0 0 35 41 2
276 33
276 114
1 1 2 0 0 0 0 13 15 0 0 3
229 70
230 70
230 60
0 2 17 0 0 0 0 0 15 35 0 3
231 33
230 33
230 42
2 1 17 0 0 8320 0 31 33 0 0 3
193 32
193 33
304 33
1 1 2 0 0 0 0 14 31 0 0 4
82 53
98 53
98 32
157 32
9 1 13 0 0 0 0 16 32 0 0 5
379 142
402 142
402 116
404 116
404 101
2 2 15 0 0 4224 0 33 32 0 0 5
340 33
403 33
403 52
404 52
404 65
2 10 18 0 0 8320 0 34 16 0 0 4
346 75
381 75
381 133
379 133
1 1 19 0 0 8320 0 34 16 0 0 4
310 75
288 75
288 133
315 133
2 2 17 0 0 0 0 35 16 0 0 3
254 114
315 114
315 142
2 3 16 0 0 4224 0 17 16 0 0 4
183 121
282 121
282 151
315 151
2 1 2 0 0 0 0 20 18 0 0 3
109 299
190 299
190 335
2 1 2 0 0 0 0 21 19 0 0 3
107 197
150 197
150 205
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
8 72 199 96
15 78 191 94
22 NAME: SHAHRIYAR SHAHID
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
516 53 627 77
523 58 619 74
12 DEMODULATION
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-05 2e-07 2e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
